`include "parameter.v" 
module VC_allocator(
    input clk,
    input rst,
    
