`include "para.v"
module reduction_tree#()
(
    input clk,
    input rst,
    input [FLIT_SIZE * N - 1 : 0] 


);
