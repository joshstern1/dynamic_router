`include "para.sv"
 module network_tb;



 	reg clk,rst;

	always #5 clk=~clk;

	network    net0(clk,rst);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_0_LOCAL.txt",net0.n_0_0_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_0_LOCAL.txt",net0.n_0_0_0.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_0_XPOS.txt",net0.n_0_0_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_0_XNEG.txt",net0.n_0_0_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_0_YPOS.txt",net0.n_0_0_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_0_YNEG.txt",net0.n_0_0_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_0_ZPOS.txt",net0.n_0_0_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_0_ZNEG.txt",net0.n_0_0_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_0_LOCAL.txt",net0.n_0_0_0.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_0_XPOS.txt",net0.n_0_0_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_0_XNEG.txt",net0.n_0_0_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_0_YPOS.txt",net0.n_0_0_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_0_YNEG.txt",net0.n_0_0_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_0_ZPOS.txt",net0.n_0_0_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_0_ZNEG.txt",net0.n_0_0_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_0_LOCAL.txt",net0.n_0_0_0.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_0_XPOS.txt",net0.n_0_0_0.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_0_XNEG.txt",net0.n_0_0_0.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_0_YPOS.txt",net0.n_0_0_0.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_0_YNEG.txt",net0.n_0_0_0.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_0_ZPOS.txt",net0.n_0_0_0.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_0_ZNEG.txt",net0.n_0_0_0.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_0_0_0.txt",net0.n_0_0_0.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_1_LOCAL.txt",net0.n_0_0_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_1_LOCAL.txt",net0.n_0_0_1.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_1_XPOS.txt",net0.n_0_0_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_1_XNEG.txt",net0.n_0_0_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_1_YPOS.txt",net0.n_0_0_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_1_YNEG.txt",net0.n_0_0_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_1_ZPOS.txt",net0.n_0_0_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_1_ZNEG.txt",net0.n_0_0_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_1_LOCAL.txt",net0.n_0_0_1.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_1_XPOS.txt",net0.n_0_0_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_1_XNEG.txt",net0.n_0_0_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_1_YPOS.txt",net0.n_0_0_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_1_YNEG.txt",net0.n_0_0_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_1_ZPOS.txt",net0.n_0_0_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_1_ZNEG.txt",net0.n_0_0_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_1_LOCAL.txt",net0.n_0_0_1.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_1_XPOS.txt",net0.n_0_0_1.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_1_XNEG.txt",net0.n_0_0_1.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_1_YPOS.txt",net0.n_0_0_1.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_1_YNEG.txt",net0.n_0_0_1.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_1_ZPOS.txt",net0.n_0_0_1.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_1_ZNEG.txt",net0.n_0_0_1.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_0_0_1.txt",net0.n_0_0_1.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_0_LOCAL.txt",net0.n_0_1_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_0_LOCAL.txt",net0.n_0_1_0.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_0_XPOS.txt",net0.n_0_1_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_0_XNEG.txt",net0.n_0_1_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_0_YPOS.txt",net0.n_0_1_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_0_YNEG.txt",net0.n_0_1_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_0_ZPOS.txt",net0.n_0_1_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_0_ZNEG.txt",net0.n_0_1_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_0_LOCAL.txt",net0.n_0_1_0.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_0_XPOS.txt",net0.n_0_1_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_0_XNEG.txt",net0.n_0_1_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_0_YPOS.txt",net0.n_0_1_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_0_YNEG.txt",net0.n_0_1_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_0_ZPOS.txt",net0.n_0_1_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_0_ZNEG.txt",net0.n_0_1_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_0_LOCAL.txt",net0.n_0_1_0.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_0_XPOS.txt",net0.n_0_1_0.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_0_XNEG.txt",net0.n_0_1_0.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_0_YPOS.txt",net0.n_0_1_0.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_0_YNEG.txt",net0.n_0_1_0.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_0_ZPOS.txt",net0.n_0_1_0.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_0_ZNEG.txt",net0.n_0_1_0.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_0_1_0.txt",net0.n_0_1_0.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_1_LOCAL.txt",net0.n_0_1_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_1_LOCAL.txt",net0.n_0_1_1.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_1_XPOS.txt",net0.n_0_1_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_1_XNEG.txt",net0.n_0_1_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_1_YPOS.txt",net0.n_0_1_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_1_YNEG.txt",net0.n_0_1_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_1_ZPOS.txt",net0.n_0_1_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_1_ZNEG.txt",net0.n_0_1_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_1_LOCAL.txt",net0.n_0_1_1.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_1_XPOS.txt",net0.n_0_1_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_1_XNEG.txt",net0.n_0_1_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_1_YPOS.txt",net0.n_0_1_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_1_YNEG.txt",net0.n_0_1_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_1_ZPOS.txt",net0.n_0_1_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_1_ZNEG.txt",net0.n_0_1_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_1_LOCAL.txt",net0.n_0_1_1.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_1_XPOS.txt",net0.n_0_1_1.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_1_XNEG.txt",net0.n_0_1_1.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_1_YPOS.txt",net0.n_0_1_1.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_1_YNEG.txt",net0.n_0_1_1.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_1_ZPOS.txt",net0.n_0_1_1.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_1_ZNEG.txt",net0.n_0_1_1.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_0_1_1.txt",net0.n_0_1_1.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_0_LOCAL.txt",net0.n_1_0_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_0_LOCAL.txt",net0.n_1_0_0.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_0_XPOS.txt",net0.n_1_0_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_0_XNEG.txt",net0.n_1_0_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_0_YPOS.txt",net0.n_1_0_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_0_YNEG.txt",net0.n_1_0_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_0_ZPOS.txt",net0.n_1_0_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_0_ZNEG.txt",net0.n_1_0_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_0_LOCAL.txt",net0.n_1_0_0.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_0_XPOS.txt",net0.n_1_0_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_0_XNEG.txt",net0.n_1_0_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_0_YPOS.txt",net0.n_1_0_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_0_YNEG.txt",net0.n_1_0_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_0_ZPOS.txt",net0.n_1_0_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_0_ZNEG.txt",net0.n_1_0_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_0_LOCAL.txt",net0.n_1_0_0.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_0_XPOS.txt",net0.n_1_0_0.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_0_XNEG.txt",net0.n_1_0_0.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_0_YPOS.txt",net0.n_1_0_0.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_0_YNEG.txt",net0.n_1_0_0.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_0_ZPOS.txt",net0.n_1_0_0.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_0_ZNEG.txt",net0.n_1_0_0.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_1_0_0.txt",net0.n_1_0_0.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_1_LOCAL.txt",net0.n_1_0_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_1_LOCAL.txt",net0.n_1_0_1.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_1_XPOS.txt",net0.n_1_0_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_1_XNEG.txt",net0.n_1_0_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_1_YPOS.txt",net0.n_1_0_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_1_YNEG.txt",net0.n_1_0_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_1_ZPOS.txt",net0.n_1_0_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_1_ZNEG.txt",net0.n_1_0_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_1_LOCAL.txt",net0.n_1_0_1.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_1_XPOS.txt",net0.n_1_0_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_1_XNEG.txt",net0.n_1_0_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_1_YPOS.txt",net0.n_1_0_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_1_YNEG.txt",net0.n_1_0_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_1_ZPOS.txt",net0.n_1_0_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_1_ZNEG.txt",net0.n_1_0_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_1_LOCAL.txt",net0.n_1_0_1.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_1_XPOS.txt",net0.n_1_0_1.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_1_XNEG.txt",net0.n_1_0_1.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_1_YPOS.txt",net0.n_1_0_1.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_1_YNEG.txt",net0.n_1_0_1.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_1_ZPOS.txt",net0.n_1_0_1.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_1_ZNEG.txt",net0.n_1_0_1.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_1_0_1.txt",net0.n_1_0_1.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_0_LOCAL.txt",net0.n_1_1_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_0_LOCAL.txt",net0.n_1_1_0.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_0_XPOS.txt",net0.n_1_1_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_0_XNEG.txt",net0.n_1_1_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_0_YPOS.txt",net0.n_1_1_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_0_YNEG.txt",net0.n_1_1_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_0_ZPOS.txt",net0.n_1_1_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_0_ZNEG.txt",net0.n_1_1_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_0_LOCAL.txt",net0.n_1_1_0.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_0_XPOS.txt",net0.n_1_1_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_0_XNEG.txt",net0.n_1_1_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_0_YPOS.txt",net0.n_1_1_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_0_YNEG.txt",net0.n_1_1_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_0_ZPOS.txt",net0.n_1_1_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_0_ZNEG.txt",net0.n_1_1_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_0_LOCAL.txt",net0.n_1_1_0.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_0_XPOS.txt",net0.n_1_1_0.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_0_XNEG.txt",net0.n_1_1_0.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_0_YPOS.txt",net0.n_1_1_0.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_0_YNEG.txt",net0.n_1_1_0.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_0_ZPOS.txt",net0.n_1_1_0.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_0_ZNEG.txt",net0.n_1_1_0.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_1_1_0.txt",net0.n_1_1_0.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_1_LOCAL.txt",net0.n_1_1_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_1_LOCAL.txt",net0.n_1_1_1.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_1_XPOS.txt",net0.n_1_1_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_1_XNEG.txt",net0.n_1_1_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_1_YPOS.txt",net0.n_1_1_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_1_YNEG.txt",net0.n_1_1_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_1_ZPOS.txt",net0.n_1_1_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_1_ZNEG.txt",net0.n_1_1_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_1_LOCAL.txt",net0.n_1_1_1.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_1_XPOS.txt",net0.n_1_1_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_1_XNEG.txt",net0.n_1_1_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_1_YPOS.txt",net0.n_1_1_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_1_YNEG.txt",net0.n_1_1_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_1_ZPOS.txt",net0.n_1_1_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_1_ZNEG.txt",net0.n_1_1_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_1_LOCAL.txt",net0.n_1_1_1.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_1_XPOS.txt",net0.n_1_1_1.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_1_XNEG.txt",net0.n_1_1_1.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_1_YPOS.txt",net0.n_1_1_1.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_1_YNEG.txt",net0.n_1_1_1.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_1_ZPOS.txt",net0.n_1_1_1.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_1_ZNEG.txt",net0.n_1_1_1.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_1_1_1.txt",net0.n_1_1_1.local_unit_inst.data);
	initial begin
		clk=0;
		rst=1;

		#100 rst=0;
	end
endmodule
