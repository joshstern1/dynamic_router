module reduction_tree#()
(
    input clk,
    input rst,
    input [FLIT_SIZE - 1 : 0] 


);
