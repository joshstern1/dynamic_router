`include "para.v"
module switch#()
(
    input clk,
    input rst,
    
);
